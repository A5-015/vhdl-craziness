----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:56:38 05/05/2019 
-- Design Name: 
-- Module Name:    display_and_controller_unit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.common.all

entity display_and_controller_unit is
Port (data_in : in STD_LOGIC_VECTOR ((instruction_width - 1) downto 0;	-- data from ROM
); 				

end display_and_controller_unit;

architecture Behavioral of display_and_controller_unit is

begin


end Behavioral;

